/*/////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
 /////////////////////////////////////////////////// SHIFT UNIT ////////////////////////////////////////////////////////////////
 //////////////////////////////////////// Developed By: Willian Analdo Nunes ///////////////////////////////////////////////////
 //////////////////////////////////////////// PUCRS, Porto Alegre, 2020      ///////////////////////////////////////////////////
 /////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////*/

//`include "pkg.sv"
import my_pkg::*;

module shiftUnit(
    input logic clk,
    input logic [31:0]  opA,
    input logic [4:0]  opB,
    input instruction_type i,
    output logic [31:0] result_out);

    logic [31:0] result;

    always_comb 
        if(i==OP0)                  // Shift logic left (SLL)
            result <= opA << opB[4:0];
        else if(i==OP1)
            result <= opA >> opB[4:0];  // Shift logic right (SRL)
        else 
            result <= $signed(opA) >>> opB[4:0]; // Shift arithmetic right (SRA)

    always @(posedge clk)
        result_out <= result;


endmodule
