/*!\file testbench.sv
 * PUCRS-RV VERSION - 1.0 - Public Release
 *
 * Distribution:  December 2021
 *
 * Willian Nunes   <willian.nunes@edu.pucrs.br>
 * Marcos Sartori  <marcos.sartori@acad.pucrs.br>
 * Ney calazans    <ney.calazans@pucrs.br>
 *
 * Research group: GAPH-PUCRS  <>
 *
 * \brief
 * Testbench for pucrs-rv simulation.
 *
 * \detailed
 * Testbench for pucrs-rv simulation.
 */

`timescale 1ns/1ps

import my_pkg::*;

///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
/////////////////////////////////////////////////////// CPU TESTBENCH IMPLEMENTATION //////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
module Testbench_With_BRAMs ();

logic         clk=1, rstCPU;
logic         enable;
logic [31:0]  data_read, DATA_address, data_write;
logic [3:0]   write;
logic [31:0]  IRQ;
byte          char;

assign IRQ = '0;
/////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
////////////////////////////////////////////////////// RESET CPU ////////////////////////////////////////////////////////////////////////////////////
/////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
    initial begin
        rstCPU = 0;
        #100 rstCPU = 1;
    end

/////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
////////////////////////////////////////////////////// Clock generator //////////////////////////////////////////////////////////////////////////////
/////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
    always begin
        #5.0 clk = 0;
        #5.0 clk = 1;
    end

/////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
////////////////////////////////////////////////////// CPU INSTANTIATION ////////////////////////////////////////////////////////////////////////////
/////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
    PUCR5_With_BRAMs dut (
        .clk(clk), 
        .reset(rstCPU), 
        .DATA_in(data_read), 
        .DATA_out(data_write), 
        .DATA_address(DATA_address),
        .enable(enable),
        .write(write),
        .IRQ(IRQ)
    );

/////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
////////////////////////////////////////////////////// Memory Mapped regs ///////////////////////////////////////////////////////////////////////////
/////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
    always @(posedge clk) 
        if(enable) begin
            ///////////////////////////////////// OUTPUT REG ///////////////////////////////////
            if((DATA_address == 32'h80004000 || DATA_address == 32'h80001000) && write!=0) begin
                char <= data_write[7:0];
                $write("%c",char);
            end
            ///////////////////////////////////// END REG //////////////////////////////////////
            if(DATA_address==32'h80000000 && write!=0) begin
                $display("# %t END OF SIMULATION",$time);
                $finish;
            end
            ///////////////////////////////////// TIMER REG ////////////////////////////////////
            if(DATA_address==32'h80006000 && write==0)
                data_read <= $time/1000;
        
        end else
            data_read <= '0;

endmodule
