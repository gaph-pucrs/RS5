import my_pkg::*;

module Peripherals (
    input logic         clk,
    input logic         reset,
    input logic         enable,
    input logic [3:0]   write,
    input logic [31:0]  DATA_address,
    input logic [31:0]  DATA_in,
    output logic [31:0] DATA_out,
    output logic [7:0]  gpioa_out,
    output logic [7:0]  gpioa_addr,
    input logic         BTND,
    output logic        UART_TX,
    output logic        stall,
    output logic [31:0] IRQ,
    input logic         Interrupt_ACK
);

logic stall_r;
logic [31:0] DATA_r, counter;
logic Buffer_write, Buffer_read, Buffer_empty, Buffer_full;
logic [7:0] Buffer_data;
logic UART_send, UART_ready;
logic [7:0] UART_data;
logic BTND_Debounced, BTND_Debounced_r, Button_Detected, Button_request;
/////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
////////////////////////////////////////////////////// Writes in Peripherals ////////////////////////////////////////////////////////////////////////
/////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
    always @(posedge clk)
        if (enable==1 && write!=0) begin
            ///////////////////////////////////// OUTPUT REG ///////////////////////////////////
            if ((DATA_address == 32'h80004000 || DATA_address == 32'h80001000) && Buffer_full==0) begin
                gpioa_out <= DATA_in[7:0];
                gpioa_addr <= 8'h84;
                Buffer_write <= 1;
                Buffer_data <= DATA_in[7:0];
            end
            ///////////////////////////////////// END REG //////////////////////////////////////
            else if (DATA_address==32'h80000000)
                gpioa_addr <= 8'h80;
            ///////////////////////////////////// NOTHING //////////////////////////////////////
            else begin
                gpioa_out <= '0;
                gpioa_addr <= '0;
                Buffer_write <= '0;         
            end

        end else begin
            gpioa_out <= '0;
            gpioa_addr <= '0;
            Buffer_write <= '0;         
        end

/////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
////////////////////////////////////////////////////// Reads from Peripherals ///////////////////////////////////////////////////////////////////////
/////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
    always @(posedge clk)
        if (enable==1 && write==0) begin
        ///////////////////////////////////// TIMER REG ////////////////////////////////////
            if (DATA_address==32'h80006000)
                DATA_r <= counter;
            else
                DATA_r <= '0;

        end else begin
            DATA_r <= '0;
        end

/////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
////////////////////////////////////////////////////// INTERRUPT CONTROL ////////////////////////////////////////////////////////////////////////////
/////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
    always @(posedge clk)
        if (reset)
            IRQ <= '0;
        ///////////////////////////////////// EXTERNAL /////////////////////////////////////
        else if (IRQ[11]==1 && Interrupt_ACK)
            IRQ[11] <= 0;
        else if (Button_request==1)
            IRQ[11] <= 1;
        ///////////////////////////////////// TIMER ////////////////////////////////////////
        else if (IRQ[7]==1 && Interrupt_ACK)
            IRQ[7] <= 0;
        else if (counter>=32'h0EE6B280)              // 1 SEC = (02FAF080)50000000 * 20ns                * 5 =  h0EE6B280
            IRQ[7] <= 1;

/////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
////////////////////////////////////////////////////// TIMER AND BUTTON /////////////////////////////////////////////////////////////////////////////
/////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
    always @(posedge clk)
        if (reset)
            counter <= 0;
        else if (IRQ[7]==1 && Interrupt_ACK)
            counter <= 0;
        else
            counter <= counter + 1;

    always @(posedge clk )
        if (reset)
            Button_request <= 0;
        else if (IRQ[11]==1 && Interrupt_ACK)
            Button_request <= 0;
        else if (Button_Detected==1 || Button_request)
            Button_request <= 1;

    debouncer #(.DEBNC_CLOCKS(2**16), .PORT_WIDTH(1)) Debouncer (
        .CLK_I(clk),
        .SIGNAL_I(BTND),
        .SIGNAL_O(BTND_Debounced)
    );

    always @(posedge clk )
        BTND_Debounced_r <= BTND_Debounced;

    assign Button_Detected = (BTND_Debounced_r==0 && BTND_Debounced==1);
/////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
////////////////////////////////////////////////////// STALL GENERATION /////////////////////////////////////////////////////////////////////////////
/////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
    always_comb
        if(enable==1) begin
            ///////////////////////////////////// READS ////////////////////////////////////////////
            if (write==0 && stall_r!=1)
                if (DATA_address==32'h80006000)
                    stall <= 1;
                else
                    stall <= 0;
            ///////////////////////////////////// WRITES ///////////////////////////////////////////
            else if (write!=0)
                if ((DATA_address == 32'h80004000 || DATA_address == 32'h80001000) && Buffer_full==1)
                    stall <= 1;
                else
                    stall <= 0;

            else
                stall <= 0;

        end else
                stall <= 0;

    always @(posedge clk) begin
        stall_r <= stall;
        DATA_out <= DATA_r;
    end

/////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
////////////////////////////////////////////////////// UART INSTANTIATION ///////////////////////////////////////////////////////////////////////////
/////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
    UART_TX_CTRL UART(
        .CLK(clk),
        .SEND(UART_send),
        .DATA(UART_data),
        .READY(UART_ready),
        .UART_TX(UART_TX)
    );

/////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
////////////////////////////////////////////////////// UART BUFFER //////////////////////////////////////////////////////////////////////////////////
/////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
    FIFO_BUFFER_UART FIFO_BUFFER_UART1 (
    .clk(clk),                // input wire clk
    .srst(reset),             // input wire srst
    .din(Buffer_data),        // input wire [7 : 0] din
    .wr_en(Buffer_write),     // input wire wr_en
    .rd_en(Buffer_read),      // input wire rd_en
    .dout(UART_data),         // output wire [7 : 0] dout
    .full(Buffer_full),       // output wire full
    .empty(Buffer_empty)      // output wire empty
    );

    assign Buffer_read = UART_ready & !Buffer_empty & !UART_send;

    always @(posedge clk ) begin
        UART_send <= Buffer_read;
    end

endmodule
