module atomic (
    input logic clk,
    input logic reset_n,
    input iTypeAtomic_e atomic_operation_i,

    output logic hold_o
);






endmodule