/*!\file testbench.sv
 * PUCRS-RV VERSION - 1.0 - Public Release
 *
 * Distribution:  December 2021
 *
 * Willian Nunes   <willian.nunes@edu.pucrs.br>
 * Marcos Sartori  <marcos.sartori@acad.pucrs.br>
 * Ney calazans    <ney.calazans@pucrs.br>
 *
 * Research group: GAPH-PUCRS  <>
 *
 * \brief
 * Testbench for pucrs-rv simulation.
 *
 * \detailed
 * Testbench for pucrs-rv simulation.
 */

`timescale 1ns/1ps

`include "../rtl/pkg.sv"
`include "../rtl/xus.sv"
`include "../rtl/fetch.sv"
`include "../rtl/decoder.sv"
`include "../rtl/execute.sv"
`include "../rtl/retire.sv"
`include "../rtl/regbank.sv"
`include "../rtl/CSRBank.sv"
`include "../rtl/PUCRS-RV.sv"
`include "./ram.sv"

import my_pkg::*;

///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
/////////////////////////////////////////////////////// CPU TESTBENCH IMPLEMENTATION //////////////////////////////////////////////////////////
///////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
module PUCRS_RV_tb ();

logic         clk=1, rstCPU;
logic [31:0]  i_address, instruction;
logic         enable_ram, enable_tb;
logic [31:0]  DATA_address, data_read, data_write;
logic [3:0]   write;
byte          char;
logic [31:0]  data_ram, data_tb;
logic [31:0]  IRQ;

////////////////////////////////////////////////////// Clock generator //////////////////////////////////////////////////////////////////////////////
    always begin
        #5.0 clk = 0;
        #5.0 clk = 1;
    end

/////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
////////////////////////////////////////////////////// CPU INSTANTIATION ////////////////////////////////////////////////////////////////////////////
/////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
    PUCRS_RV dut (
        .clk(clk), 
        .reset(rstCPU), 
        .instruction(instruction), 
        .i_address(i_address), 
        .enable(enable_int), 
        .write(write),
        .DATA_address(DATA_address),
        .DATA_in(data_read), 
        .DATA_out(data_write),
        .IRQ(IRQ)
    );

/////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
////////////////////////////////////////////////////// RAM INSTANTIATION ///////////////////////////////////////////////////////////////////////
/////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
    RAM_mem RAM_MEM(
        .clk(clk), 
        .rst(rstCPU), 
        .en(enable_ram), 
        .i_data(instruction),
        .w_en(write), 
        .i_addr(i_address[15:0]), 
        .d_addr(DATA_address[15:0]), 
        .w_data(data_write), 
        .r_data(data_ram)
    );

    assign enable_tb = (DATA_address > 32'h0000FFFF && enable_int) ? 1 : 0;
    assign enable_ram = (DATA_address <= 32'h0000FFFF && enable_int) ? 1 : 0;

    assign data_read = (enable_tb) ? data_tb : data_ram;

/////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
////////////////////////////////////////////////////// Memory Mapped regs ///////////////////////////////////////////////////////////////////////////
/////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
    always @(posedge clk)
        if(enable_tb) begin
            ///////////////////////////////////// OUTPUT REG ///////////////////////////////////
            if((DATA_address == 32'h80004000 || DATA_address == 32'h80001000) && write!=0) begin
                char <= data_write[7:0];
                $write("%c",char);
            end
            ///////////////////////////////////// END REG //////////////////////////////////////
            if(DATA_address==32'h80000000 && write!=0) begin
                $display("# %t END OF SIMULATION",$time);
                $finish;
            end
            ///////////////////////////////////// TIMER REG ////////////////////////////////////
            if(DATA_address==32'h80006000 && write==0)
                data_tb <= $time/1000;
        
        end else
                data_tb <= '0;

/////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
////////////////////////////////////////////////////// TIMER generator //////////////////////////////////////////////////////////////////////////////
/////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
integer TIMER;
    always @(posedge clk or negedge rstCPU) begin
        if (!rstCPU)
            TIMER <= 0;
        else begin
            TIMER <= TIMER + 1;
//            if(TIMER % 500 == 0)
//                IRQ[7] <= 1;
        end
    end

/////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
////////////////////////////////////////////////////// RESET CPU ////////////////////////////////////////////////////////////////////////////////////
/////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
    initial begin
        rstCPU = 0;                                          // RESET for CPU initialization
        IRQ <= '0;
        
        #100 rstCPU = 1;                                     // Hold state for 100 ns
/*
        #300
        IRQ[11] <= 1;
        #70
        IRQ[11] <= 0;
        #30
        IRQ[3] <= 1;
        #70
        IRQ[3] <= 0;
        #30
        IRQ[7] <= 1;
        #70
        IRQ[7] <= 0;
        #70
        IRQ[7] <= 'Z;
*/
    end

endmodule
