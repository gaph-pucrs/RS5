`timescale 1ns/1ns

`include "../rtl/RS5_pkg.sv"

module tb_top
    import RS5_pkg::*;
;

    logic        clk=1, reset_n;

    testbench #(
        .INSTRUCTION_SET(RV32M),
        .USE_XOSVM(1'b1),
        .USE_ZIHPM(1'b1)
    ) tb (
        .clk_i(clk),
        .reset_n(reset_n)
    );

///////////////////////////////////////// Clock generator //////////////////////////////
    always begin
        #5.0 clk = 0;
        #5.0 clk = 1;
    end

/////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
////////////////////////////////////////////////////// RESET CPU ////////////////////////////////////////////////////////////////////////////////////
/////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
    initial begin
        reset_n = 0;                                          // RESET for CPU initialization

        #100 reset_n = 1;                                     // Hold state for 100 ns
    end

endmodule
